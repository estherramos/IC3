library IEEE;
use IEEE.std_logic_1164.all;

Entity ejercicio1_a is
    port(
        x,y,z: in std_logic;
        F1: out std_logic;
	    F2: out std_logic
    );
end entity ejercicio1_a;



